module main

import core { Vector3, Quaternion }

fn main() {
	dump(f32(1))
}
