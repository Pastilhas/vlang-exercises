module core

pub interface Component {}
