module main

import core { Vector3, Quaternion }

fn main() {
	v := Vector3.new(1,0,0)
	q := Quaternion.new(0, 0.707, 0, 0.707)

	dump(f32(1))
}
