module core

pub interface Component {
	component_id string

}
